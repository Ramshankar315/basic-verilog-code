module notgate(input A,output Y);
assign Y=!A;
endmodule
