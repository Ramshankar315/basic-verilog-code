module AND_2 (output Y, input A, B);
assign Y = A & B; 
endmodule
